module trim_gen (CLK50,RST,DOUT,TRIMCODE);
    input CLK50, RST;
    output reg DOUT;
    output reg [11:0] TRIMCODE;

    
    
endmodule